//You are given a dynamic array of integers where each element can have a value between 0 and 100. You are required to write a function in SystemVerilog that:

//Randomizes the dynamic array (with values between 0 and 100).
//Computes the sum of all the even numbers in the array using array reduction methods.
//Additionally, compute the sum of all the elements at odd indices.
